module Display(
    input           i_rst_n;
    input           i_clk;
    input [19:0]    i_addr;
    input [19:0]    i_addr_end;
);


endmodule